*** SPICE deck for cell critical_path{sch} from library Assignment4
*** Created on Mon Oct 30, 2023 15:57:41
*** Last revised on Wed Dec 06, 2023 21:24:32
*** Written on Wed Dec 06, 2023 21:24:40 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.01FF

*** SUBCIRCUIT NAND2__NAND2 FROM CELL NAND2:NAND2{sch}
.SUBCKT NAND2__NAND2 A B Y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@2 net@22 A gnd gnd nmos L=0.022U W=0.176U
Mnmos@3 Y B net@22 gnd nmos L=0.022U W=0.176U
Mpmos@2 vdd B Y vdd pmos L=0.022U W=0.176U
Mpmos@3 vdd A Y vdd pmos L=0.022U W=0.176U

* Spice Code nodes in cell cell 'NAND2:NAND2{sch}'
.include "E:\IITM Acads\Sem 5\DIC\Electric\22nm_HP.pm"
.ENDS NAND2__NAND2

*** SUBCIRCUIT Assignment3__assignment3_new FROM CELL Assignment3:assignment3_new{sch}
.SUBCKT Assignment3__assignment3_new A B Ci Co_ S_
** GLOBAL gnd
** GLOBAL vdd
Mnmos@12 Co_ Ci net@88 gnd nmos L=0.022U W=0.088U
Mnmos@13 net@88 B gnd gnd nmos L=0.022U W=0.088U
Mnmos@14 net@69 Ci gnd gnd nmos L=0.022U W=0.088U
Mnmos@15 net@69 Ci gnd gnd nmos L=0.022U W=0.088U
Mnmos@16 net@69 Ci gnd gnd nmos L=0.022U W=0.088U
Mnmos@17 net@69 B gnd gnd nmos L=0.022U W=0.088U
Mnmos@18 net@69 B gnd gnd nmos L=0.022U W=0.088U
Mnmos@19 net@69 B gnd gnd nmos L=0.022U W=0.088U
Mnmos@20 Co_ A net@69 gnd nmos L=0.022U W=0.088U
Mnmos@21 Co_ A net@69 gnd nmos L=0.022U W=0.088U
Mnmos@22 Co_ A net@69 gnd nmos L=0.022U W=0.088U
Mnmos@23 net@64 A gnd gnd nmos L=0.022U W=0.088U
Mnmos@24 net@64 B gnd gnd nmos L=0.022U W=0.088U
Mnmos@25 net@64 Ci gnd gnd nmos L=0.022U W=0.088U
Mnmos@26 S_ Co_ net@64 gnd nmos L=0.022U W=0.088U
Mnmos@27 S_ A net@60 gnd nmos L=0.022U W=0.132U
Mnmos@28 net@60 B net@142 gnd nmos L=0.022U W=0.132U
Mnmos@29 net@142 Ci gnd gnd nmos L=0.022U W=0.132U
Mpmos@12 vdd B net@108 vdd pmos L=0.022U W=0.176U
Mpmos@13 net@108 Ci Co_ vdd pmos L=0.022U W=0.176U
Mpmos@14 vdd Ci net@115 vdd pmos L=0.022U W=0.176U
Mpmos@15 vdd Ci net@115 vdd pmos L=0.022U W=0.176U
Mpmos@16 vdd Ci net@115 vdd pmos L=0.022U W=0.176U
Mpmos@17 vdd B net@115 vdd pmos L=0.022U W=0.176U
Mpmos@18 vdd B net@115 vdd pmos L=0.022U W=0.176U
Mpmos@19 vdd B net@115 vdd pmos L=0.022U W=0.176U
Mpmos@20 net@115 A Co_ vdd pmos L=0.022U W=0.176U
Mpmos@21 net@115 A Co_ vdd pmos L=0.022U W=0.176U
Mpmos@22 net@115 A Co_ vdd pmos L=0.022U W=0.176U
Mpmos@23 vdd A net@55 vdd pmos L=0.022U W=0.176U
Mpmos@24 vdd B net@55 vdd pmos L=0.022U W=0.176U
Mpmos@25 vdd Ci net@55 vdd pmos L=0.022U W=0.176U
Mpmos@26 net@55 Co_ S_ vdd pmos L=0.022U W=0.176U
Mpmos@27 vdd Ci net@61 vdd pmos L=0.022U W=0.264U
Mpmos@28 net@61 B net@63 vdd pmos L=0.022U W=0.264U
Mpmos@29 net@63 A S_ vdd pmos L=0.022U W=0.264U

* Spice Code nodes in cell cell 'Assignment3:assignment3_new{sch}'
.include "E:\IITM Acads\Sem 5\DIC\Electric\22nm_HP.pm"
*.param vdd = 0.8
*v1 vdd gnd DC {vdd}
*v2 A gnd PULSE(0 {vdd} 400p 100p 100p 400p 1n)
*v3 B gnd PULSE(0 {vdd} 900p 100p 100p 900p 2n)
*v4 Ci gnd PULSE(0 {vdd} 1900p 100p 100p 1900p 4n)
*.tran 0 8n
.ENDS Assignment3__assignment3_new

*** SUBCIRCUIT NAND2__inverter FROM CELL NAND2:inverter{sch}
.SUBCKT NAND2__inverter INP OUT
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT INP gnd gnd nmos L=0.022U W=0.088U
Mpmos@0 vdd INP OUT vdd pmos L=0.022U W=0.176U

* Spice Code nodes in cell cell 'NAND2:inverter{sch}'
.include "E:\IITM Acads\Sem 5\DIC\Electric\22nm_HP.pm"
*v1 vdd gnd DC 0.8
*v2 INP gnd pwl(0 0 100p 0.8 1n 0.8 1.1n 0 2n 0)
*.tran 2.1n
*.END
.ENDS NAND2__inverter

.global gnd vdd

*** TOP LEVEL CELL: Assignment4:critical_path{sch}
XNAND2@2 c vdd net@267 NAND2__NAND2
Xassignme@7 net@15 b1 gnd net@281 net@78 Assignment3__assignment3_new
Xassignme@8 net@281 b1 a1 net@286 assignme@8_S_ Assignment3__assignment3_new
Xassignme@9 net@286 b1 a1 net@290 net@80 Assignment3__assignment3_new
Xassignme@10 net@290 b1 a1 net@295 assignme@10_S_ Assignment3__assignment3_new
Xassignme@11 net@295 b1 a1 net@299 net@81 Assignment3__assignment3_new
Xassignme@12 net@299 b1 a1 net@302 assignme@12_S_ Assignment3__assignment3_new
Xassignme@13 net@302 b1 a1 net@306 net@83 Assignment3__assignment3_new
Xassignme@14 net@306 b1 a1 co s Assignment3__assignment3_new
Xassignme@15 c1 gnd a1 net@137 net@134 Assignment3__assignment3_new
Xassignme@16 net@134 b net@188 net@317 net@119 Assignment3__assignment3_new
Xassignme@17 net@119 b net@218 net@140 net@107 Assignment3__assignment3_new
Xassignme@18 net@107 b net@195 net@142 net@126 Assignment3__assignment3_new
Xassignme@19 net@126 b net@230 net@144 net@110 Assignment3__assignment3_new
Xassignme@20 net@110 b net@233 net@146 net@111 Assignment3__assignment3_new
Xassignme@21 net@111 b net@209 net@148 net@15 Assignment3__assignment3_new
Xassignme@22 a b net@137 assignme@22_Co_ assignme@22_S_ Assignment3__assignment3_new
Xassignme@23 a b net@317 assignme@23_Co_ assignme@23_S_ Assignment3__assignment3_new
Xassignme@24 a b net@140 assignme@24_Co_ assignme@24_S_ Assignment3__assignment3_new
Xassignme@25 a b net@142 assignme@25_Co_ assignme@25_S_ Assignment3__assignment3_new
Xassignme@26 a b net@144 assignme@26_Co_ assignme@26_S_ Assignment3__assignment3_new
Xassignme@27 a b net@146 assignme@27_Co_ assignme@27_S_ Assignment3__assignment3_new
Xassignme@28 a b net@148 assignme@28_Co_ assignme@28_S_ Assignment3__assignment3_new
Xinverter@3 net@78 inverter@3_OUT NAND2__inverter
Xinverter@4 net@80 inverter@4_OUT NAND2__inverter
Xinverter@5 net@81 inverter@5_OUT NAND2__inverter
Xinverter@6 net@83 inverter@6_OUT NAND2__inverter
Xinverter@8 a a1 NAND2__inverter
Xinverter@9 a net@188 NAND2__inverter
Xinverter@10 a net@218 NAND2__inverter
Xinverter@11 a net@195 NAND2__inverter
Xinverter@12 a net@230 NAND2__inverter
Xinverter@13 a net@233 NAND2__inverter
Xinverter@14 a net@209 NAND2__inverter
Xinverter@15 net@267 c1 NAND2__inverter

* Spice Code nodes in cell cell 'Assignment4:critical_path{sch}'
.include "E:\IITM Acads\Sem 5\DIC\Electric\22nm_HP.pm"
.param vdd=0.8
v1 vdd gnd DC {vdd}
v2 a1 gnd DC 0
v3 b1 gnd DC {vdd}
v4 a gnd DC {vdd}
v5 b gnd DC {vdd}
v6 c gnd PULSE(0 {vdd} 900p 100p 100p 900p 2n)
.meas tran cr
+trig v(c) = {vdd}/2 cross =1
+targ v(s) = {vdd}/2 cross =1
.meas tran cf
+trig v(c) = {vdd}/2 cross =2
+targ v(s) = {vdd}/2 cross =2
.tran 0 4n
